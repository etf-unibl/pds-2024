
library ieee;
use ieee.std_logic_1164.all;

entity test is
	port
	(
		i1	: in  std_logic;
		o1	: out std_logic
	);
end test;

architecture test_arch of test is
begin
	
end test_arch;