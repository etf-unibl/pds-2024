library ieee;
use ieee.std_logic_1164.all;

entity invertor is
	port
	(
		input	: in  std_logic;
		output	: out std_logic
	);
end invertor;

architecture in_arch of invertor is
begin
	
end in_arch;