library ieee;
use ieee.std_logic_1164.all;

entity test is
	port
	(
		test_input	: in  std_logic;
		test_output	: out std_logic
	);
end test;

architecture test_arch of test is
begin
end test_arch;